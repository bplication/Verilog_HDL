module DOT(S,B,clk, dot_14, dot_10);

input clk;
input [2:0] S;
input [2:0] B;
output [13:0] dot_14;
output [9:0] dot_10;
reg [13:0] dot_14;
reg [9:0] dot_10;
reg [3:0] count_10;
reg CLK0;
reg [7:0] CLK_COUNT0;
reg state;
reg [3:0] h_state;
reg [31:0] dot_count;
reg dot_clk;
reg [4:0] dot_state;

initial
begin 
 	dot_10 <= 10'b1000000000;
	dot_14 <= 14'b00000000000000;
end

parameter SS = 0;
parameter BB = 1;
	
always @(negedge clk) // CLK/0
	if (CLK_COUNT0==100) begin CLK_COUNT0<=0; CLK0<=1; end
	else begin CLK_COUNT0 <= CLK_COUNT0+1; CLK0<=0; end
	
	
	always@(posedge CLK0)
		if(count_10 >= 10) count_10 <= 0;
		else count_10 <= count_10 + 1;
	
	always@(posedge CLK0)
		state <= !state;

	always@(posedge clk)
		if (dot_count==2500000) begin dot_count<=0; dot_clk<=1; end
		else begin dot_count <= dot_count+1; dot_clk<=0; end
		
	always@(posedge dot_clk)
		h_state <= h_state+1;


	always@(count_10) //��� seg ���� 
		case(count_10)
		1:  dot_10 <= 10'b1000000000; //line1
		2:  dot_10 <= 10'b0100000000; //line2
		3:  dot_10 <= 10'b0010000000; //line3
		4:  dot_10 <= 10'b0001000000;  //line4
		5:  dot_10 <= 10'b0000100000;  //line5
		6:  dot_10 <= 10'b0000010000;  //line6
		7:  dot_10 <= 10'b0000001000;  //line7
		8:  dot_10 <= 10'b0000000100;  //line8
		9:  dot_10 <= 10'b0000000010;  //line9
		10:  dot_10 <= 10'b0000000001; //line1
		endcase
	
//1,2��и�,����,S
always@(*)
	begin
	if(S<4)
	begin
	case(state)
	SS : case(S)

		0 : case (count_10)
			1: dot_14 <= 14'b00000000000000;
			2: dot_14 <= 14'b11111110000000;
			3: dot_14 <= 14'b10000010000000;
			4: dot_14 <= 14'b11111110000000;
			5: dot_14 <= 14'b00000000000000;
			6: dot_14 <= 14'b11110010000000; //s line6
			7: dot_14 <= 14'b10010010000000; //s line7
			8: dot_14 <= 14'b10010010000000; //s line8
			9: dot_14 <= 14'b10010010000000; //s line9
			10: dot_14 <= 14'b10011110000000; //s line10
			endcase
		
		1 : case (count_10)
			1: dot_14 <= 14'b00100010000000;
			2: dot_14 <= 14'b01000010000000;
			3: dot_14 <= 14'b11111110000000;
			4: dot_14 <= 14'b00000010000000;
			5: dot_14 <= 14'b00000010000000;
			6: dot_14 <= 14'b11110010000000; //s line6
			7: dot_14 <= 14'b10010010000000; //s line7
			8: dot_14 <= 14'b10010010000000; //s line8
			9: dot_14 <= 14'b10010010000000; //s line9
			10: dot_14 <= 14'b10011110000000; //s line10
			endcase
		
		2 : case(count_10)
			1: dot_14 <= 14'b10011110000000; //line1
			2: dot_14 <= 14'b10010010000000; //line2
			3: dot_14 <= 14'b10010010000000; //line3
			4: dot_14 <= 14'b10010010000000; //line4
 			5: dot_14 <= 14'b11110010000000; //line5
			6: dot_14 <= 14'b11110010000000; //s line6
			7: dot_14 <= 14'b10010010000000; //s line7
			8: dot_14 <= 14'b10010010000000; //s line8
			9: dot_14 <= 14'b10010010000000; //s line9
			10: dot_14 <= 14'b10011110000000; //s line10
			endcase

		3 : case(count_10)
			1: dot_14 <= 14'b10010010000000; //line1
			2: dot_14 <= 14'b10010010000000; //line2
			3: dot_14 <= 14'b10010010000000; //line3	
			4: dot_14 <= 14'b10010010000000; //line4		
			5: dot_14 <= 14'b11111110000000; //line5		
			6: dot_14 <= 14'b11110010000000; //s line6
			7: dot_14 <= 14'b10010010000000; //s line7
			8: dot_14 <= 14'b10010010000000; //s line8
			9: dot_14 <= 14'b10010010000000; //s line9
			10: dot_14 <= 14'b10011110000000; //s line10
			endcase

		4 : case(count_10)
			1: dot_14 <= 14'b11110000000000; //4 line1
			2: dot_14 <= 14'b00010000000000; //4 line2
			3: dot_14 <= 14'b00010000000000; //4 line3
			4: dot_14 <= 14'b00010000000000; //4 line4
			5: dot_14 <= 14'b11111110000000; //4 line5
			6: dot_14 <= 14'b11110010000000; //s line6
			7: dot_14 <= 14'b10010010000000; //s line7 
			8: dot_14 <= 14'b10010010000000; //s line8
			9: dot_14 <= 14'b10010010000000; //s line9
			10: dot_14 <= 14'b10011110000000; //s line10
			endcase
		
		default : case (count_10)
			1: dot_14 <= 14'b00000000000000;
			2: dot_14 <= 14'b00000000000000;
			3: dot_14 <= 14'b00000000000000;
			4: dot_14 <= 14'b00000000000000;
			5: dot_14 <= 14'b00000000000000;
			6: dot_14 <= 14'b11110010000000; //s line6
			7: dot_14 <= 14'b10010010000000; //s line7
			8: dot_14 <= 14'b10010010000000; //s line8
			9: dot_14 <= 14'b10010010000000; //s line9
			10: dot_14 <= 14'b10011110000000; //s line10
			endcase
		endcase
	
	BB : case(B)
	
		0 : case (count_10)
			1: dot_14 <= 14'b00000000000000;
			2: dot_14 <= 14'b00000001111111;
			3: dot_14 <= 14'b00000001000001;
			4: dot_14 <= 14'b00000001111111;
			5: dot_14 <= 14'b00000000000000;
			6: dot_14 <= 14'b00000001111111; //B line6
			7: dot_14 <= 14'b00000001001001; //B line7
			8: dot_14 <= 14'b00000001001001; //B line8
			9: dot_14 <= 14'b00000001001001; //B line9
			10: dot_14 <= 14'b00000000110110; //B line10
			endcase
			
		1 : case(count_10)
			1: dot_14 <= 14'b00000000010001; //line1
			2: dot_14 <= 14'b00000000100001; //line2
			3: dot_14 <= 14'b00000001111111; //line3
			4: dot_14 <= 14'b00000000000001; //line4
			5: dot_14 <= 14'b00000000000001; //line5
			6: dot_14 <= 14'b00000001111111; //B line6
			7: dot_14 <= 14'b00000001001001; //B line7
			8: dot_14 <= 14'b00000001001001; //B line8
			9: dot_14 <= 14'b00000001001001; //B line9
			10: dot_14 <= 14'b00000000110110; //B line10
			endcase
	
		2 : case(count_10)
			1: dot_14 <= 14'b00000001001111; //line1
			2: dot_14 <= 14'b00000001001001; //line2
			3: dot_14 <= 14'b00000001001001; //line3
			4: dot_14 <= 14'b00000001001001; //line4
			5: dot_14 <= 14'b00000001111001; //line5
			6: dot_14 <= 14'b00000001111111; //B line6
			7: dot_14 <= 14'b00000001001001; //B line7
			8: dot_14 <= 14'b00000001001001; //B line8
			9: dot_14 <= 14'b00000001001001; //B line9
			10: dot_14 <= 14'b00000000110110; //B line10
			endcase

	
		3 : case(count_10)
			1: dot_14 <= 14'b00000001001001; //line1
			2: dot_14 <= 14'b00000001001001; //line2
			3: dot_14 <= 14'b00000001001001; //line3
			4: dot_14 <= 14'b00000001001001; //line4
			5: dot_14 <= 14'b00000001111111; //line5
			6: dot_14 <= 14'b00000001111111; //B line6
			7: dot_14 <= 14'b00000001001001; //B line7
			8: dot_14 <= 14'b00000001001001; //B line8
			9: dot_14 <= 14'b00000001001001; //B line9
			10: dot_14 <= 14'b00000000110110; //B line10
			endcase

		4 : case(count_10)		
			1: dot_14 <= 14'b00000001111000; //line1
			2: dot_14 <= 14'b00000000001000; //line2
			3: dot_14 <= 14'b00000000001000; //line3
			4: dot_14 <= 14'b00000000001000; //line4
			5: dot_14 <= 14'b00000001111111; //line5
			6: dot_14 <= 14'b00000001111111; //B line6
			7: dot_14 <= 14'b00000001001001; //B line7
			8: dot_14 <= 14'b00000001001001; //B line8
			9: dot_14 <= 14'b00000001001001; //B line9
			10: dot_14 <= 14'b00000000110110; //B line10
			endcase

		default : case (count_10)
			1: dot_14 <= 14'b00000000000000;
			2: dot_14 <= 14'b00000000000000;
			3: dot_14 <= 14'b00000000000000;
			4: dot_14 <= 14'b00000000000000;
			5: dot_14 <= 14'b00000000000000;
			6: dot_14 <= 14'b00000001111111; //B line6
			7: dot_14 <= 14'b00000001001001; //B line7
			8: dot_14 <= 14'b00000001001001; //B line8
			9: dot_14 <= 14'b00000001001001; //B line9
			10: dot_14 <= 14'b00000000110110; //B line10
			endcase
			
		endcase
	endcase
	end
	
	else if(S==4)
	begin	
	case(h_state)
	0: case(count_10)
		1: dot_14 <= 14'b00000000000000;
		2: dot_14 <= 14'b00000000000000;
		3: dot_14 <= 14'b00000000000000;
		4: dot_14 <= 14'b00000111100000;
		5: dot_14 <= 14'b00000111100000;
		6: dot_14 <= 14'b00000111100000;
		7: dot_14 <= 14'b00000111100000;
		8: dot_14 <= 14'b00000000000000;
		9: dot_14 <= 14'b00000000000000;
		10: dot_14 <= 14'b00000000000000;
		endcase

	1: case(count_10)
		1: dot_14 <= 14'b00000000000000;
		2: dot_14 <= 14'b00000000000000;
		3: dot_14 <= 14'b00000000000000;
		4: dot_14 <= 14'b00000111100000;
		5: dot_14 <= 14'b00001100110000;
		6: dot_14 <= 14'b00001100110000;
		7: dot_14 <= 14'b00000111100000;
		8: dot_14 <= 14'b00000000000000;
		9: dot_14 <= 14'b00000000000000;
		10: dot_14 <= 14'b00000000000000;
		endcase

	2: case(count_10)
		1: dot_14 <= 14'b00000000000000;
		2: dot_14 <= 14'b00011111111000;
		3: dot_14 <= 14'b00110000001100;
		4: dot_14 <= 14'b01100000000110;
		5: dot_14 <= 14'b01100000000110;
		6: dot_14 <= 14'b01100000000110;
		7: dot_14 <= 14'b01100000000110;
		8: dot_14 <= 14'b00110000001100;
		9: dot_14 <= 14'b00011111111000;
		10: dot_14 <= 14'b00000000000000;
		endcase

	3: case(count_10)
		1: dot_14 <= 14'b00111111111100;
		2: dot_14 <= 14'b01100000000110;
		3: dot_14 <= 14'b11000000000011;
		4: dot_14 <= 14'b11000000000011;
		5: dot_14 <= 14'b11000000000011;
		6: dot_14 <= 14'b11000000000011;
		7: dot_14 <= 14'b11000000000011;
		8: dot_14 <= 14'b11000000000011;
		9: dot_14 <= 14'b01100000000110;
		10: dot_14 <= 14'b00111111111100;
		endcase

	4: case(count_10)
		1: dot_14 <= 14'b00001110000000;
		2: dot_14 <= 14'b00010000001110;
		3: dot_14 <= 14'b00001000010000;
		4: dot_14 <= 14'b00000100100000;
		5: dot_14 <= 14'b00000011000000;
		6: dot_14 <= 14'b00000011000000;
		7: dot_14 <= 14'b00000100100000;
		8: dot_14 <= 14'b00001000010000;
		9: dot_14 <= 14'b11110000001000;
		10: dot_14 <= 14'b00000001110000;
		endcase

	5: case(count_10)
		1: dot_14 <= 14'b00000111000000;
		2: dot_14 <= 14'b00001000001110;
		3: dot_14 <= 14'b00000100010001;
		4: dot_14 <= 14'b00000100100001;
		5: dot_14 <= 14'b00000011000001;
		6: dot_14 <= 14'b00000111000000;
		7: dot_14 <= 14'b10001001000000;
		8: dot_14 <= 14'b10010000100000;
		9: dot_14 <= 14'b11100000010000;
		10: dot_14 <= 14'b00000111100000;
		endcase


	6: case(count_10)
		1: dot_14 <= 14'b00000011110000;
		2: dot_14 <= 14'b00000010000000;
		3: dot_14 <= 14'b10000010000000;
		4: dot_14 <= 14'b10000010000000;
		5: dot_14 <= 14'b10000011111111;
		6: dot_14 <= 14'b11111111000001;
		7: dot_14 <= 14'b00000001000001;
		8: dot_14 <= 14'b00000001000001;
		9: dot_14 <= 14'b00000001000000;
		10: dot_14 <= 14'b00001111000000;
		endcase


	7: case(count_10)
		1: dot_14 <= 14'b00111100011110;
		2: dot_14 <= 14'b01000000100000;
		3: dot_14 <= 14'b00100001000000;
		4: dot_14 <= 14'b00011100100000;
		5: dot_14 <= 14'b00000011000000;
		6: dot_14 <= 14'b00000011000000;
		7: dot_14 <= 14'b10001100110000;
		8: dot_14 <= 14'b10010000001000;
		9: dot_14 <= 14'b10100000000100;
		10: dot_14 <= 14'b11000000011110;
		endcase


	8: case(count_10)
		1: dot_14 <= 14'b00000011110000;
		2: dot_14 <= 14'b00000010000000;
		3: dot_14 <= 14'b10000010000000;
		4: dot_14 <= 14'b10000010000000;
		5: dot_14 <= 14'b10000011111111;
		6: dot_14 <= 14'b11111111000001;
		7: dot_14 <= 14'b00000001000001;
		8: dot_14 <= 14'b00000001000001;
		9: dot_14 <= 14'b00000001000000;
		10: dot_14 <= 14'b00001111000000;
		endcase


	9: case(count_10)
		1: dot_14 <= 14'b00000111000000;
		2: dot_14 <= 14'b00001000001110;
		3: dot_14 <= 14'b00000100010001;
		4: dot_14 <= 14'b00000100100001;
		5: dot_14 <= 14'b00000011000001;
		6: dot_14 <= 14'b00000111000000;
		7: dot_14 <= 14'b10001001000000;
		8: dot_14 <= 14'b10010000100000;
		9: dot_14 <= 14'b11100000010000;
		10: dot_14 <= 14'b00000111100000;
		endcase


	10: case(count_10)
		1: dot_14 <= 14'b00001110000000;
		2: dot_14 <= 14'b00010000001110;
		3: dot_14 <= 14'b00001000010000;
		4: dot_14 <= 14'b00000100100000;
		5: dot_14 <= 14'b00000011000000;
		6: dot_14 <= 14'b00000011000000;
		7: dot_14 <= 14'b00000100100000;
		8: dot_14 <= 14'b00001000010000;
		9: dot_14 <= 14'b11110000001000;
		10: dot_14 <= 14'b00000001110000;
		endcase

	11: case(count_10)
		1: dot_14 <= 14'b00001110000000;
		2: dot_14 <= 14'b00010000001110;
		3: dot_14 <= 14'b00001000010000;
		4: dot_14 <= 14'b00000100100000;
		5: dot_14 <= 14'b00000011000000;
		6: dot_14 <= 14'b00000011000000;
		7: dot_14 <= 14'b00000100100000;
		8: dot_14 <= 14'b00001000010000;
		9: dot_14 <= 14'b11110000001000;
		10: dot_14 <= 14'b00000001110000;
		endcase
		
	12: case(count_10)
		1: dot_14 <= 14'b00000111000000;
		2: dot_14 <= 14'b00001000001110;
		3: dot_14 <= 14'b00000100010001;
		4: dot_14 <= 14'b00000100100001;
		5: dot_14 <= 14'b00000011000001;
		6: dot_14 <= 14'b00000111000000;
		7: dot_14 <= 14'b10001001000000;
		8: dot_14 <= 14'b10010000100000;
		9: dot_14 <= 14'b11100000010000;
		10: dot_14 <= 14'b00000111100000;
		endcase

	13: case(count_10)
		1: dot_14 <= 14'b00000011110000;
		2: dot_14 <= 14'b00000010000000;
		3: dot_14 <= 14'b10000010000000;
		4: dot_14 <= 14'b10000010000000;
		5: dot_14 <= 14'b10000011111111;
		6: dot_14 <= 14'b11111111000001;
		7: dot_14 <= 14'b00000001000001;
		8: dot_14 <= 14'b00000001000001;
		9: dot_14 <= 14'b00000001000000;
		10: dot_14 <= 14'b00001111000000;
		endcase

	14: case(count_10)
		1: dot_14 <= 14'b00111100011110;
		2: dot_14 <= 14'b01000000100000;
		3: dot_14 <= 14'b00100001000000;
		4: dot_14 <= 14'b00011100100000;
		5: dot_14 <= 14'b00000011000000;
		6: dot_14 <= 14'b00000011000000;
		7: dot_14 <= 14'b10001100110000;
		8: dot_14 <= 14'b10010000001000;
		9: dot_14 <= 14'b10100000000100;
		10: dot_14 <= 14'b11000000011110;
		endcase

	15: case(count_10)
		1: dot_14 <= 14'b11000000000011;
		2: dot_14 <= 14'b11000000000011;
		3: dot_14 <= 14'b11000000000011;
		4: dot_14 <= 14'b11000000000011;
		5: dot_14 <= 14'b11111111111111;
		6: dot_14 <= 14'b11111111111111;
		7: dot_14 <= 14'b11000000000011;
		8: dot_14 <= 14'b11000000000011;
		9: dot_14 <= 14'b11000000000011;
		10: dot_14 <= 14'b11000000000011;
		endcase
	endcase
	end
	end


endmodule